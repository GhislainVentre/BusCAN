LIBRARY ieee;
  USE ieee.std_logic_1164.ALL;
  USE ieee.numeric_std.ALL;

Entity Transmitter is
port(
	clk	: in std_logic;
	Tx		: out std_logic
);
end entity;

architecture Behavioral of Transmitter is
begin
end architecture;
