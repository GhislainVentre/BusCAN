library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity Gestionnaire_de_protocole_CAN is
end entity;

architecture arc of Gestionnaire_de_protocole_CAN is
begin

end architecture;